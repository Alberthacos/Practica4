NET"' LOC="";
NET"' LOC="";